library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Full_Adder is
	port
	(
		A	:	in	std_logic;
		B	:	in	std_logic;
		Cin	:	in	std_logic;
		Sum	:	out	std_logic;
		Cout	:	out	std_logic
	);
end Full_Adder;


architecture behaviour of Full_Adder is
begin
	process(A, B, Cin)
	begin
		Sum 	<= (A xor B xor Cin);
		Cout 	<= (A and B) or (B and Cin) or (A and Cin);
	end process;
end behaviour;
