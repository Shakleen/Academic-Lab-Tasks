library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Or_Gate is
	port
	(
		A, B	:	in	std_logic;
		C	:	out	std_logic
	);
end Or_Gate;


architecture behaviour of Or_Gate is
begin
	process(A, B)
	begin
		C <= A or B;
	end process;
end behaviour;